module s1_2class_easy_hybrid2_seed22(
  input  wire [112:0] in_bits,
  output wire [1:0] out_bits
);

  wire input_1 = in_bits[0];
  wire input_2 = in_bits[1];
  wire input_3 = in_bits[2];
  wire input_4 = in_bits[3];
  wire input_5 = in_bits[4];
  wire input_6 = in_bits[5];
  wire input_7 = in_bits[6];
  wire input_8 = in_bits[7];
  wire input_9 = in_bits[8];
  wire input_10 = in_bits[9];
  wire input_11 = in_bits[10];
  wire input_12 = in_bits[11];
  wire input_13 = in_bits[12];
  wire input_14 = in_bits[13];
  wire input_15 = in_bits[14];
  wire input_16 = in_bits[15];
  wire input_17 = in_bits[16];
  wire input_18 = in_bits[17];
  wire input_19 = in_bits[18];
  wire input_20 = in_bits[19];
  wire input_21 = in_bits[20];
  wire input_22 = in_bits[21];
  wire input_23 = in_bits[22];
  wire input_24 = in_bits[23];
  wire input_25 = in_bits[24];
  wire input_26 = in_bits[25];
  wire input_27 = in_bits[26];
  wire input_28 = in_bits[27];
  wire input_29 = in_bits[28];
  wire input_30 = in_bits[29];
  wire input_31 = in_bits[30];
  wire input_32 = in_bits[31];
  wire input_33 = in_bits[32];
  wire input_34 = in_bits[33];
  wire input_35 = in_bits[34];
  wire input_36 = in_bits[35];
  wire input_37 = in_bits[36];
  wire input_38 = in_bits[37];
  wire input_39 = in_bits[38];
  wire input_40 = in_bits[39];
  wire input_41 = in_bits[40];
  wire input_42 = in_bits[41];
  wire input_43 = in_bits[42];
  wire input_44 = in_bits[43];
  wire input_45 = in_bits[44];
  wire input_46 = in_bits[45];
  wire input_47 = in_bits[46];
  wire input_48 = in_bits[47];
  wire input_49 = in_bits[48];
  wire input_50 = in_bits[49];
  wire input_51 = in_bits[50];
  wire input_52 = in_bits[51];
  wire input_53 = in_bits[52];
  wire input_54 = in_bits[53];
  wire input_55 = in_bits[54];
  wire input_56 = in_bits[55];
  wire input_57 = in_bits[56];
  wire input_58 = in_bits[57];
  wire input_59 = in_bits[58];
  wire input_60 = in_bits[59];
  wire input_61 = in_bits[60];
  wire input_62 = in_bits[61];
  wire input_63 = in_bits[62];
  wire input_64 = in_bits[63];
  wire input_65 = in_bits[64];
  wire input_66 = in_bits[65];
  wire input_67 = in_bits[66];
  wire input_68 = in_bits[67];
  wire input_69 = in_bits[68];
  wire input_70 = in_bits[69];
  wire input_71 = in_bits[70];
  wire input_72 = in_bits[71];
  wire input_73 = in_bits[72];
  wire input_74 = in_bits[73];
  wire input_75 = in_bits[74];
  wire input_76 = in_bits[75];
  wire input_77 = in_bits[76];
  wire input_78 = in_bits[77];
  wire input_79 = in_bits[78];
  wire input_80 = in_bits[79];
  wire input_81 = in_bits[80];
  wire input_82 = in_bits[81];
  wire input_83 = in_bits[82];
  wire input_84 = in_bits[83];
  wire input_85 = in_bits[84];
  wire input_86 = in_bits[85];
  wire input_87 = in_bits[86];
  wire input_88 = in_bits[87];
  wire input_89 = in_bits[88];
  wire input_90 = in_bits[89];
  wire input_91 = in_bits[90];
  wire input_92 = in_bits[91];
  wire input_93 = in_bits[92];
  wire input_94 = in_bits[93];
  wire input_95 = in_bits[94];
  wire input_96 = in_bits[95];
  wire input_97 = in_bits[96];
  wire input_98 = in_bits[97];
  wire input_99 = in_bits[98];
  wire input_100 = in_bits[99];
  wire input_101 = in_bits[100];
  wire input_102 = in_bits[101];
  wire input_103 = in_bits[102];
  wire input_104 = in_bits[103];
  wire input_105 = in_bits[104];
  wire input_106 = in_bits[105];
  wire input_107 = in_bits[106];
  wire input_108 = in_bits[107];
  wire input_109 = in_bits[108];
  wire input_110 = in_bits[109];
  wire input_111 = in_bits[110];
  wire input_112 = in_bits[111];
  wire input_113 = in_bits[112];
  wire const_114 = 1'b1;
  wire const_115 = 1'b0;

  wire gate_l1_116 = (input_82 | input_17);
  wire gate_l1_117 = (input_1 & input_2 & input_3);
  wire gate_l1_118 = 1'b1;
  wire gate_l1_119 = (((input_36 ? 1 : 0)) >= 1);
  wire gate_l1_120 = (input_24 ^ input_84);
  wire gate_l1_121 = (((input_1 ? 1 : 0) + (input_2 ? 1 : 0)) >= 1);
  wire gate_l1_122 = (((input_1 ? 1 : 0)) >= 1);
  wire gate_l1_123 = ((input_16 & input_65) | (input_16 & (1'b0)));
  wire gate_l1_124 = (((input_1 ? 1 : 0) + (input_2 ? 1 : 0)) >= 1);
  wire gate_l1_125 = 1'b1;
  wire gate_l1_126 = (input_1 | input_2);
  wire gate_l1_127 = (input_1 | (input_2 & (input_3 | input_4 | input_5 | input_6 | input_7 | input_8 | input_9 | input_10 | input_11 | input_12 | input_13 | input_14 | input_15 | input_16 | input_17 | input_18 | input_19 | input_20 | input_21 | input_22 | input_23 | input_24 | input_25 | input_26 | input_27 | input_28 | input_29 | input_30 | input_31 | input_32 | input_33 | input_34 | input_35 | input_36 | input_37 | input_38 | input_39 | input_40 | input_41 | input_42 | input_43 | input_44 | input_45 | input_46 | input_47 | input_48 | input_49 | input_50 | input_51 | input_52 | input_53 | input_54 | input_55 | input_56 | input_57 | input_58 | input_59 | input_60 | input_61 | input_62 | input_63 | input_64 | input_65 | input_66 | input_67 | input_68 | input_69 | input_70 | input_71 | input_72 | input_73 | input_74 | input_75 | input_76 | input_77 | input_78 | input_79 | input_80 | input_81 | input_82 | input_83 | input_84 | input_85 | input_86 | input_87 | input_88 | input_89 | input_90 | input_91 | input_92 | input_93 | input_94 | input_95 | input_96 | input_97 | input_98 | input_99 | input_100 | input_101 | input_102 | input_103 | input_104 | input_105 | input_106 | input_107 | input_108 | input_109 | input_110 | input_111 | input_112 | input_113 | const_114 | const_115)));
  wire gate_l1_128 = (((input_1 ? 1 : 0) + (input_2 ? 1 : 0)) >= 1);
  wire gate_l1_129 = 1'b0;
  wire gate_l1_130 = (input_90 & input_9);
  wire gate_l1_131 = (input_1 | (input_2 & (input_3 | input_4 | input_5 | input_6 | input_7 | input_8 | input_9 | input_10 | input_11 | input_12 | input_13 | input_14 | input_15 | input_16 | input_17 | input_18 | input_19 | input_20 | input_21 | input_22 | input_23 | input_24 | input_25 | input_26 | input_27 | input_28 | input_29 | input_30 | input_31 | input_32 | input_33 | input_34 | input_35 | input_36 | input_37 | input_38 | input_39 | input_40 | input_41 | input_42 | input_43 | input_44 | input_45 | input_46 | input_47 | input_48 | input_49 | input_50 | input_51 | input_52 | input_53 | input_54 | input_55 | input_56 | input_57 | input_58 | input_59 | input_60 | input_61 | input_62 | input_63 | input_64 | input_65 | input_66 | input_67 | input_68 | input_69 | input_70 | input_71 | input_72 | input_73 | input_74 | input_75 | input_76 | input_77 | input_78 | input_79 | input_80 | input_81 | input_82 | input_83 | input_84 | input_85 | input_86 | input_87 | input_88 | input_89 | input_90 | input_91 | input_92 | input_93 | input_94 | input_95 | input_96 | input_97 | input_98 | input_99 | input_100 | input_101 | input_102 | input_103 | input_104 | input_105 | input_106 | input_107 | input_108 | input_109 | input_110 | input_111 | input_112 | input_113 | const_114 | const_115)));
  wire gate_l1_132 = (((input_1 ? 1 : 0) + (input_2 ? 1 : 0) + (input_3 ? 1 : 0) + (input_4 ? 1 : 0)) >= 2);
  wire gate_l1_133 = (((input_54 ? 1 : 0) + (input_27 ? 1 : 0) + (input_107 ? 1 : 0) + (input_87 ? 1 : 0)) >= 2);
  wire gate_l1_134 = (input_15 | (input_5 & (input_97)));
  wire gate_l1_135 = 1'b0;
  wire gate_l1_136 = (input_67 ^ input_11);
  wire gate_l1_137 = (input_68 ^ input_81);
  wire gate_l1_138 = (((input_56 ? 1 : 0) + (input_28 ? 1 : 0)) >= 1);
  wire gate_l1_139 = (input_1 & input_2);
  wire gate_l2_140 = (((input_85 ? 1 : 0) + (input_107 ? 1 : 0) + (input_60 ? 1 : 0) + (input_92 ? 1 : 0)) >= 2);
  wire gate_l2_141 = 1'b1;
  wire gate_l2_142 = (input_95 & input_57);
  wire gate_l2_143 = (gate_l1_119 | input_28);
  wire gate_l2_144 = (input_84 ^ gate_l1_124);
  wire gate_l2_145 = (((input_1 ? 1 : 0) + (input_2 ? 1 : 0)) >= 1);
  wire gate_l2_146 = (input_81 | input_10);
  wire gate_l2_147 = (input_96 & input_111);
  wire gate_l2_148 = (((input_56 ? 1 : 0) + (gate_l1_136 ? 1 : 0)) >= 1);
  wire gate_l2_149 = (gate_l1_122 & input_79);
  wire gate_l2_150 = ((input_7 & input_28) | (input_7 & (input_50 | input_42)));
  wire gate_l2_151 = (input_49 & input_99);
  wire output_0_152 = (((input_108 ? 1 : 0) + (input_91 ? 1 : 0)) >= 1);
  wire output_1_153 = 1'b1;

  assign out_bits[0] = output_0_152;
  assign out_bits[1] = output_1_153;
endmodule
